module matrix_mac_unit;

endmodule
