module matrix_mac_unit(
    clock,
    reset
    );

endmodule