//===========================================//
//  Copyright (c) Aleksandar Kostovic 2018   //
//    Matrix Multiply and Accumulate unit    //
//===========================================//

module matrix_mac_unit #(
    parameter DATA_WIDTH = 8
)( //ports
    clock,         //|<input
    reset,         //|<input
    enable,        //|<input
    clear          //|<input
);
//inputs

//outputs

//regs and/or wires

//sequential logic

//combinational logic


endmodule
