//===========================================
// Copyright (c) Aleksandar Kostovic 2018 
//   Matrix Multiply and Accumulate unit     
//===========================================

module matrix_mac_unit #(
    parameter DATA_WITDH = 8
)( //ports
    clock,         //|<input
    reset          //|<input
);

endmodule
