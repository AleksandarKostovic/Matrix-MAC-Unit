//===========================================
// Copyright (c) Aleksandar Kostovic 2018 
//   Matrix Multiply and Accumulate unit     
//===========================================

module matrix_mac_unit #(
    parameter integer DATA_WITDH = 8
)( //ports
    i_clk,       //|<i
    i_rst        //|<i
);

endmodule
