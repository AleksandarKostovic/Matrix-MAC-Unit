//===========================================
// Copyright (c) Aleksandar Kostovic 2018 
//   Matrix Multiply and Accumulate unit     
//===========================================

module matrix_mac_unit(
    clk                 //|<input
   ,rst                 //|<input
    );

endmodule
